// Verilog test fixture created from schematic /home/lamd/Documents/csse232/1516a-csse232-frenchkt-knightcm-lamd-peterseo/cla/cla.sch - Thu Nov  5 11:35:07 2015

`timescale 1ns / 1ps

module cla_cla_sch_tb();

// Inputs

// Output

// Bidirs

// Instantiate the UUT
   cla UUT (
		
   );
// Initialize Inputs
   `ifdef auto_init
       initial begin
   `endif
endmodule
